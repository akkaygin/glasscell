`default_nettype none

module glasscell(
  input Clock,
  input Reset


);

endmodule